package apb_pkg;

   import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_transaction.svh"
  `include "apb_sequencer.svh"

  `include "monitor_apb.svh"
  `include "driver_apb.svh"
  `include "agent_apb.svh"
  `include "apb_seq_lib.svh"

endpackage