package mem_pkg;

   import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "mem_transaction.svh"
  //`include "memory_coverage.svh"

  `include "mem_driver_a.svh"
  `include "mem_driver_b.svh"
  `include "mem_driver_c.svh"

  `include "mem_monitor_a.svh"
  `include "mem_monitor_b.svh"
  `include "mem_monitor_c.svh"
  `include "mem_agent.svh"

endpackage


