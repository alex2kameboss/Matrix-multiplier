module matrix_multiplier(
    input           clk     ,
    input           rst_n   
);

wrapper wrapper_i (
    .clk  ,
    .rst_n
);

endmodule