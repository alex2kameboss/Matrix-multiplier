package apb_pkg;

   import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_transaction.sv"

  `include "monitor_apb.sv"
  `include "driver_apb.sv"
  `include "agent_apb.sv"

endpackage