package env_pkg;

   import uvm_pkg::*;
   import apb_pkg::*;
   import mem_pkg::*;

   `include "uvm_macros.svh"

   `include "environment.svh"
endpackage