package test_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh";

import apb_pkg::*;
import mem_pkg::*; 
import env_pkg::*;

`include "tests_lib.svh";

    
endpackage : test_pkg